library ieee;
use ieee.std_logic_1164.all;

PACKAGE opcodes IS

	CONSTANT NOP  : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"00";
	CONSTANT SUBA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"01";
	CONSTANT CMPA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"02";
	CONSTANT LDAI : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"03";
	CONSTANT LDAD : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"04";
	CONSTANT LDAX : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"05";
	CONSTANT LDAF : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"06";
	CONSTANT STAD : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"07";
	CONSTANT STAX : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"08";
	CONSTANT STAF : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"09";
	CONSTANT JSR : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0A";
	CONSTANT RTS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0B";
	CONSTANT LINK : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0C";
	CONSTANT UNLINK : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0D";
	CONSTANT BEQ : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0E";
	CONSTANT BLT : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0F";
	CONSTANT BLE : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"10";
	CONSTANT BRA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"11";
	CONSTANT ADDA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"12";
	CONSTANT CLRA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"13";
	CONSTANT PUSHA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"14";
	CONSTANT PUSHX : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"15";
	CONSTANT POPA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"16";
	CONSTANT POPX : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"17";
	CONSTANT INCA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"18";
	CONSTANT DECA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"19";
	CONSTANT INCX : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1A";
	CONSTANT DECX : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1B";
	CONSTANT SHRA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1C";
	CONSTANT SHLA : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1D";
	CONSTANT HALT : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1E";
	CONSTANT SHRL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1F";
END PACKAGE;